,0
0,Alabama
1,Arizona
2,Arkansas
3,Colorado
4,Connecticut
5,Delaware
6,Georgia
7,Idaho
8,Illinois
9,Iowa
10,Kansas
11,Kentucky
12,Louisiana
13,Maine
14,Maryland
15,Massachusetts
16,Michigan
17,Minnesota
18,Mississippi
19,Missouri
20,Montana
21,Nebraska
22,Nevada
23,New Hampshire
24,New Jersey
25,New Mexico
26,New York
27,North Carolina
28,North Dakota
29,Oklahoma
30,Oregon
31,Pennsylvania
32,Rhode Island
33,South Carolina
34,South Dakota
35,Tennessee
36,Utah
37,Vermont
38,Virginia
39,Washington
40,West Virginia
41,Wisconsin
42,Wyoming
